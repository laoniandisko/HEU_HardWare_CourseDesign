library verilog;
use verilog.vl_types.all;
entity computer1119_vlg_vec_tst is
end computer1119_vlg_vec_tst;
