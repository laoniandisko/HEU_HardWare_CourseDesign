library verilog;
use verilog.vl_types.all;
entity SHEFT_vlg_vec_tst is
end SHEFT_vlg_vec_tst;
