library verilog;
use verilog.vl_types.all;
entity uControl1119_vlg_vec_tst is
end uControl1119_vlg_vec_tst;
