library verilog;
use verilog.vl_types.all;
entity move_computer1119_vlg_vec_tst is
end move_computer1119_vlg_vec_tst;
